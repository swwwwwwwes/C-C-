change for git hub
