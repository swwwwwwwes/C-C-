ahb is the advanced high performance bus

ram is using BRAM concept to implement,

//try to test the branch merge!
