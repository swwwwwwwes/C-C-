ahb is the advanced high performance bus
